/*
	Autor: Albert Espi�a Rojas
	Modulo: I2C_SLAVE_ADDRESS_MATCH

Modulo para comprovar si el slave tiene la direcci�n de memor�a la cual solicita el master.
El modulo dispone de dos funciones seleccionables con la variable modo. La primera es comprovar si el dispositivo
tiene esa direcci�n de memoria como hemos mencionado anteriormente o si queremos a�adir una nueva direcci�n de memoria.
Para ello habr� la posibilidad de tener diferentes direcciones de memoria, las cuales no tienen porque ser consecutivas
y debido a que habr� un tama�o fijado de direcciones, se proceder� a actuar como LIFO.No obstante el a�adir memorias ser� recomendable
hacerlo al inicio del programa como una configuraci�n previa.

*/

module I2C_SLAVE_ADDRESS_MATCH #( parameter LENGTH, parameter MaxAddress)(Clk, Rst, Enable, Mode, InputAddress, AddressFound);
	input Clk;
 	input Rst; 
	input Enable; 
	input Mode;
	input [LENGTH - 1: 0]InputAddress;
	output reg [LENGTH - 1: 0]AddressFound;
	reg [(LENGTH - 1)*MaxAddress: 0]AddressList;
always @(posedge Clk)
begin
    	if (!Rst) AddressFound = 1'b0;
  	else if (Enable) begin
		if (Mode) AddressFound = 1'b0; //Falta a�adir cosas
		else AddressFound = 1'b0; //Falta a�adir cosas
	end
end

endmodule